/**
 * @file cordic_sine.sv
 * @author Geeoon Chung
 * @brief this file implements the cordic_sine module
 */

module cordic_sine
    #(parameter BIT_WIDTH={},
      parameter K={})
    (clk, angle, output);
    /**
     * @brief 
     */
endmodule  // cordic_sine
